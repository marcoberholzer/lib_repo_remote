cs_component_b