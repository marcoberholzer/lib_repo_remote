cs_component_a