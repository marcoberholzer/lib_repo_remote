cl_component_b
change 1