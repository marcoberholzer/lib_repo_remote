cl_component_b