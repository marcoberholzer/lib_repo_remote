cs_component_a
change 2 (branch_1)