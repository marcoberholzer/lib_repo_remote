cl_component_a