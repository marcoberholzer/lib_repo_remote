cl_component_a
change 3